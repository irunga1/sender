<?xml version="1.0" encoding="UTF-8" standalone="no"?>
<!-- Created with Inkscape (http://www.inkscape.org/) -->
<svg
    xmlns:inkscape="http://www.inkscape.org/namespaces/inkscape"
    xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"
    xmlns="http://www.w3.org/2000/svg"
    xmlns:xlink="http://www.w3.org/1999/xlink"
    xmlns:ns1="http://sozi.baierouge.fr"
    xmlns:cc="http://creativecommons.org/ns#"
    xmlns:dc="http://purl.org/dc/elements/1.1/"
    xmlns:sodipodi="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd"
    id="svg2"
    sodipodi:docname="he-man.svg"
    viewBox="0 0 153.68 258.51"
    version="1.1"
    inkscape:version="0.48.4 r9939"
  >
  <title
      id="title3003"
    >he-man</title
  >
  <sodipodi:namedview
      id="base"
      bordercolor="#666666"
      inkscape:pageshadow="2"
      inkscape:window-y="-8"
      fit-margin-left="0"
      pagecolor="#ffffff"
      inkscape:window-height="706"
      inkscape:window-maximized="1"
      inkscape:zoom="2.8"
      inkscape:window-x="-8"
      showgrid="false"
      borderopacity="1.0"
      inkscape:current-layer="layer1"
      inkscape:cx="58.286879"
      inkscape:cy="163.64145"
      fit-margin-top="0"
      fit-margin-right="0"
      fit-margin-bottom="0"
      inkscape:window-width="1366"
      inkscape:pageopacity="0.0"
      inkscape:document-units="px"
  />
  <g
      id="layer1"
      inkscape:label="Layer 1"
      inkscape:groupmode="layer"
      transform="translate(259.7 20.762)"
    >
    <path
        id="path3001"
        sodipodi:nodetypes="ccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccc"
        style="stroke-linejoin:round;fill-rule:evenodd;stroke:#d05244;stroke-width:2;fill:#090a14"
        inkscape:connector-curvature="0"
        d="m-191.93-18.232c-7.6303-0.63376-10.22 9.0204-17.076 10.154-1.8248 1.7079 0.81385 6.1632-3.0525 5.5871-1.6399 1.1473 1.7662 2.2483 0.27541 3.8715-0.39224 1.9772 0.72325 3.8199 2.2492 4.3584 0.0708 2.8964-3.9898 8.0822-6.3804 3.9875-1.6668-1.3528-1.9065-5.0628-4.7509-3.8252-3.0312-0.53011-4.2137-3.7696-4.8427-6.213-3.1169 1.4915-1.2216 6.4304 0.16885 8.7649 0.73174 2.9105 5.5495 6.6932 2.9755 9.6887-5.5936 3.4702-12.746 1.7194-16.938-3.1297-1.6387-1.5303-5.0847-2.8433-5.2788 0.60276-1.311 7.5859-0.60002 15.444 0.75739 22.882-2.231 5.6077-2.1489 12.035-5.7837 17.179-5.032 6.0129-3.936 14.56-4.3378 21.908 0.33732 5.4753 3.6474 10.201 3.9476 15.741 0.71778 2.7012 3.3055 4.8992 1.291 7.8935-1.0194 1.5597-3.7087-3.1701-6.1796-2.0283-4.2191 0.76963-2.0856 7.6044 1.8361 6.6071 3.9764 0.7858 8.5109 3.4172 7.4591 8.2299 1.3625 4.3808 7.5773 3.9588 10.695 6.4217 0.87613 2.3031-4.149 2.7856-2.341 5.5407 2.378 4.7418 8.4072 3.7474 12.738 4.3584 0.87507 7.0283-0.53476 15.074-5.2099 20.47-5.3903 3.3312-10.447 7.3847-13.587 12.959-3.4961 2.4124-8.9527 5.7046-6.5411 10.803 0.59902 6.7366 8.0679 10.12 7.8493 17.132-0.0199 6.7123 2.0169 14.498-2.3869 20.239-1.166 3.9119-3.6552 7.0577-7.3903 8.74-4.8564 3.3513-2.882 10.503 1.9279 12.82 2.5931 2.3214 5.832 2.2482 8.5837 0.20863 4.8469-2.3117 11.555-5.1018 10.594-11.771 1.1487-7.7088 0.71301-15.577 1.8687-23.235 1.5113-6.6159 5.7626-11.881 11.085-15.834 4.9141-3.4616 4.7448-9.9298 2.2951-14.837-2.8456-6.3079 4.0844-10.62 6.3345-15.764 4.27-3.7625 7.0063-8.762 9.7772-13.608 7.6064 1.3384 14.677 4.9642 21.758 7.9054 0.56228 5.2449 1.4319 11.019-2.349 15.342-2.5716 5.7722-10.612 10.253-7.4971 17.461 2.3972 2.1188 4.0209 5.4054 7.023 7.1403 5.489 5.4385 1.1241 13.35 1.4526 19.933-0.30564 4.196-0.57603 8.3946-0.85588 12.592 4.3772 3.3042 10.444 2.2667 14.299 6.4448 5.7784 3.704 13.675 4.3575 20.036 2.2256 1.1111-3.1465-3.8148-5.1771-5.5181-7.2254-4.3159-3.8124-7.9706-8.4726-11.672-12.758-0.44354-1.6679-2.957-2.0985-2.823-4.4279-2.2352-6.9341 0.13326-14.484 5.646-19.126 5.3013-3.3379 7.3879-11.041 3.259-16.112-1.1744-3.2841-3.1632-7.2142-2.4558-10.595 16.816 7.1298 32.07 18.835 50.309 22.163 0.97759-1.5789-2.5658-3.4782-3.3968-4.7293-13.838-12.231-31.302-19.198-46.132-29.929-2.4915-5.2773 2.3328-11.004 2.0426-16.506 0.71556-4.7414-0.84455-10.217 1.0099-14.559 3.239-0.25452 4.576 5.4501 8.2624 3.0833 4.7908-0.65015 7.3672-2.9662 5.9296-8.0676 0.13241-10.414-0.37409-20.906-2.5099-31.065 0.82057-6.7325-2.6762-12.603-6.6329-17.642-1.1204-3.3188 0.70309-7.2653-1.8131-10.34-2.3996-6.3894-1.5221-15.011-8.4001-18.825-3.8937-3.3994-9.9981-2.1323-12.922-6.8621-2.1771-3.6079-8.394-3.0903-8.3313-8.1836 1.3104-4.6167 8.2214-6.9835 6.9312-12.774-1.8329-7.0449-3.8751-14.987-9.387-20.03-2.3401-1.4684-5.2284-1.4882-7.8952-1.4373zm-32.407 81.836c2.8933 0.84096 2.8652 5.0302 5.8984 5.4712 1.9349 3.5856 7.1996 4.6979 8.8458 7.8543 0.36469 7.0935-6.4988 11.633-6.39 18.644-0.62615 2.7303-2.0522 5.6302-4.2689 6.9549 1.7168 3.999-5.451 2.4723-4.7738-0.6723-0.29364-1.2835 2.4958-2.2155-0.18361-2.0865-3.119-0.70598-3.7518 5.309-6.2657 1.6692-4.1816-3.6037-2.0193-10.171-2.4558-14.999 0.55521-4.748 4.6619-8.9077 2.4099-13.979-0.98873-2.1984-2.9383-6.0032 1.1246-6.1435 2.2056-0.45168 3.9689-2.1513 6.0591-2.7124zm58.342 5.2625c4.3706 3.4089-0.43222 9.9723 2.3181 14.327 3.4652 5.2583 9.6661 8.9095 10.374 15.695 1.9682 2.2122 1.1267 4.6267-0.64263 6.6303-1.2916 2.1894-1.5597 6.7535-2.1359 7.1487-2.245-7.1224-5.4152-14.013-7.1593-21.267-4.145-5.7781-9.8215-13.011-7.2296-20.563 1.6848-1.9413 1.8376-5.383 4.4755-1.9705z"
    />
  </g
  >
  <metadata
    >
    <rdf:RDF
      >
      <cc:Work
        >
        <dc:format
          >image/svg+xml</dc:format
        >
        <dc:type
            rdf:resource="http://purl.org/dc/dcmitype/StillImage"
        />
        <cc:license
            rdf:resource="http://creativecommons.org/licenses/publicdomain/"
        />
        <dc:publisher
          >
          <cc:Agent
              rdf:about="http://openclipart.org/"
            >
            <dc:title
              >Openclipart</dc:title
            >
          </cc:Agent
          >
        </dc:publisher
        >
      </cc:Work
      >
      <cc:License
          rdf:about="http://creativecommons.org/licenses/publicdomain/"
        >
        <cc:permits
            rdf:resource="http://creativecommons.org/ns#Reproduction"
        />
        <cc:permits
            rdf:resource="http://creativecommons.org/ns#Distribution"
        />
        <cc:permits
            rdf:resource="http://creativecommons.org/ns#DerivativeWorks"
        />
      </cc:License
      >
    </rdf:RDF
    >
  </metadata
  >
</svg
>
